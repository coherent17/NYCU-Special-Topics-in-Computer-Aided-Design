
module           c17 (N1, N2, N3,N6, 
    N7 , N22, 

    N23);

   wire  n8,n9
//
,
 n10,
n11 , n12
;
	input               N1, N2,N3
 , N6,N7;

	output /*fdsg*//*htrghr*/ N22,
	 	N/*;*/23;
    /*
        Hello
        // World!
    */
// gthytjthgj juythjuhyfj

    /*
        Hello
        // World!*/
    NOR2X1
U8 (./*(fdfsgsku*/A1(n8),   .A2(n9),  .ZN(N23));
	  NOR2X1 U9 /*ffffgfg/*ddasdda*/(.A1(N2), /*stshrsrhadas*/.A2(N7), .ZN(n9));//dhjikb/*
	INVX1 U10 (.I(n10), /*AAAAdsadsadsad*/ .ZN(n8));   //dghsrthrsu/*hstrtsrhrsgg?*/
    // dasdsadsadsad
            NANDX1 U11 (.A1(n11), .A2(n12),
             .ZN(N22)); //dsadsadsdsadsad
	NANDX1                   U12 (.A1(N2),   /*aaas
    dsad*/ .A2(n10), .ZN(n12))/*
      ggg
            NANDX1 U11 (.A1(n11), .A2(n12),
/*
  */;   //dshshshrshshf*/
	    /*asdhtrshbsbshsa*/NANDX1 U13 (.A1(N6),
          .A2(N3), .ZN(n10));
	NANDX1              U14    ( .A1(N1), .A2(N3), /*sagtrshyrjhrd*/.ZN(n11));
endmodule